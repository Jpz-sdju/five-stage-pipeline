module mem_wb (
    
);
    
endmodule