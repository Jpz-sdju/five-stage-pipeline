`include "para.v"
module ysyx_22040384_tiny_adder (
    input [`ysyx_22040383_width] a,
    input [`ysyx_22040383_width] b,
    output [`ysyx_22040383_width] c
);
    assign c = a+b;    
endmodule