`include "para.v"
module wb (
    input [`width] wri
);
    
endmodule