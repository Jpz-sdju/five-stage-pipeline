`include "para.v"
module ex_mem (
    input ex_is_write_dmem,
    input [1:0]ex_wb_selece,
    input [7:0] ex_write_width,
    input [`width] ex_dmem_write_data,
    input ex_pc_sel
);
    
endmodule